module tb;

$display("hi");
endmodule
